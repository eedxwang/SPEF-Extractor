module secc ( gnd, vdd, in1, in5, in9, in13, in17, in21, in25, in29, in33, in37, in41, in45, in49, in53, in57, in61, in65, in69, in73, in77, in81, in85, in89, in93, in97, in101, in105, in109, in113, in117, in121, in125, in129, in130, in131, in132, in133, in134, in135, in136, in137, out724, out725, out726, out727, out728, out729, out730, out731, out732, out733, out734, out735, out736, out737, out738, out739, out740, out741, out742, out743, out744, out745, out746, out747, out748, out749, out750, out751, out752, out753, out754, out755);

input gnd, vdd;
input in1;
input in5;
input in9;
input in13;
input in17;
input in21;
input in25;
input in29;
input in33;
input in37;
input in41;
input in45;
input in49;
input in53;
input in57;
input in61;
input in65;
input in69;
input in73;
input in77;
input in81;
input in85;
input in89;
input in93;
input in97;
input in101;
input in105;
input in109;
input in113;
input in117;
input in121;
input in125;
input in129;
input in130;
input in131;
input in132;
input in133;
input in134;
input in135;
input in136;
input in137;
output out724;
output out725;
output out726;
output out727;
output out728;
output out729;
output out730;
output out731;
output out732;
output out733;
output out734;
output out735;
output out736;
output out737;
output out738;
output out739;
output out740;
output out741;
output out742;
output out743;
output out744;
output out745;
output out746;
output out747;
output out748;
output out749;
output out750;
output out751;
output out752;
output out753;
output out754;
output out755;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_0_), .B(_538_), .Y(_412_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_535_), .C(in17), .Y(_413_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(in17), .Y(_414_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_1_), .B(_528_), .Y(_415_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_415_), .C(_545_), .Y(_416_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_416_), .Y(_4_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_548_), .C(in21), .Y(_417_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(in21), .Y(_418_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_415_), .C(_552_), .Y(_419_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_419_), .Y(_5_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_397_), .C(in25), .Y(_420_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(in25), .Y(_421_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_421_), .B(_415_), .C(_403_), .Y(_422_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_422_), .Y(_6_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_406_), .C(in29), .Y(_423_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(in29), .Y(_424_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_415_), .C(_410_), .Y(_425_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_425_), .Y(_7_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_3_), .B(_540_), .Y(_426_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_533_), .C(_426_), .Y(_427_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_427_), .C(in33), .Y(_428_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(in33), .Y(_429_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_2_), .B(_530_), .Y(_430_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_543_), .C(_430_), .Y(_431_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_539_), .C(_431_), .Y(_432_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_432_), .Y(_8_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_547_), .C(_426_), .Y(_433_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_433_), .C(in37), .Y(_434_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(in37), .Y(_435_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_551_), .C(_430_), .Y(_436_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_539_), .C(_436_), .Y(_437_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_434_), .B(_437_), .Y(_9_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_395_), .C(_426_), .Y(_438_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_438_), .C(in41), .Y(_439_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(in41), .Y(_440_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_401_), .C(_430_), .Y(_441_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_539_), .C(_441_), .Y(_442_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_442_), .Y(_10_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_405_), .C(_426_), .Y(_443_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_443_), .C(in45), .Y(_444_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(in45), .Y(_445_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_409_), .C(_430_), .Y(_446_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_445_), .B(_539_), .C(_446_), .Y(_447_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_444_), .B(_447_), .Y(_11_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_427_), .C(in49), .Y(_448_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(in49), .Y(_449_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_415_), .C(_431_), .Y(_450_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_448_), .B(_450_), .Y(_12_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_433_), .C(in53), .Y(_451_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(in53), .Y(_452_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_452_), .B(_415_), .C(_436_), .Y(_453_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_453_), .Y(_13_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_438_), .C(in57), .Y(_454_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(in57), .Y(_455_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_415_), .C(_441_), .Y(_456_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_454_), .B(_456_), .Y(_14_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_443_), .C(in61), .Y(_457_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(in61), .Y(_458_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_458_), .B(_415_), .C(_446_), .Y(_459_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_459_), .Y(_15_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_1_), .B(Ckt499b_M1_S_0_), .Y(_460_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_531_), .C(_533_), .Y(_461_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_461_), .C(in65), .Y(_462_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(in65), .Y(_463_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_1_), .B(Ckt499b_M1_S_0_), .Y(_464_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_541_), .C(_543_), .Y(_465_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_395_), .C(_465_), .Y(_466_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_466_), .Y(_16_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_533_), .C(_426_), .Y(_467_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_467_), .C(in69), .Y(_468_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(in69), .Y(_469_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_543_), .C(_430_), .Y(_470_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_469_), .B(_395_), .C(_470_), .Y(_471_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_468_), .B(_471_), .Y(_17_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_3_), .B(Ckt499b_M1_S_2_), .Y(_472_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_539_), .C(_533_), .Y(_473_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_473_), .C(in73), .Y(_474_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(in73), .Y(_475_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_3_), .B(Ckt499b_M1_S_2_), .Y(_476_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_529_), .C(_543_), .Y(_477_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_395_), .C(_477_), .Y(_478_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_478_), .Y(_18_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_533_), .C(_415_), .Y(_479_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_479_), .C(in77), .Y(_480_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(in77), .Y(_481_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_543_), .C(_412_), .Y(_482_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_481_), .B(_395_), .C(_482_), .Y(_483_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_480_), .B(_483_), .Y(_19_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_461_), .C(in81), .Y(_484_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(in81), .Y(_485_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_405_), .C(_465_), .Y(_486_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_484_), .B(_486_), .Y(_20_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_467_), .C(in85), .Y(_487_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(in85), .Y(_488_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_488_), .B(_405_), .C(_470_), .Y(_489_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_489_), .Y(_21_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_473_), .C(in89), .Y(_490_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(in89), .Y(_491_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_491_), .B(_405_), .C(_477_), .Y(_492_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_490_), .B(_492_), .Y(_22_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_479_), .C(in93), .Y(_493_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(in93), .Y(_494_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_405_), .C(_482_), .Y(_495_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_493_), .B(_495_), .Y(_23_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_531_), .C(_547_), .Y(_496_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_496_), .C(in97), .Y(_497_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(in97), .Y(_498_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_541_), .C(_551_), .Y(_499_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_395_), .C(_499_), .Y(_500_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_500_), .Y(_24_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_460_), .B(_547_), .C(_426_), .Y(_501_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_501_), .C(in101), .Y(_502_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(in101), .Y(_503_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_551_), .C(_430_), .Y(_504_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_395_), .C(_504_), .Y(_505_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_502_), .B(_505_), .Y(_25_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_539_), .C(_547_), .Y(_506_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_506_), .C(in105), .Y(_507_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(in105), .Y(_508_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_529_), .C(_551_), .Y(_509_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_395_), .C(_509_), .Y(_510_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_510_), .Y(_26_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_547_), .C(_415_), .Y(_511_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_511_), .C(in109), .Y(_512_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(in109), .Y(_513_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_551_), .C(_412_), .Y(_514_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_513_), .B(_395_), .C(_514_), .Y(_515_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_515_), .Y(_27_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_496_), .C(in113), .Y(_516_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(in113), .Y(_517_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_517_), .B(_405_), .C(_499_), .Y(_518_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_516_), .B(_518_), .Y(_28_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_501_), .C(in117), .Y(_519_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(in117), .Y(_520_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_520_), .B(_405_), .C(_504_), .Y(_521_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_521_), .Y(_29_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_506_), .C(in121), .Y(_522_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(in121), .Y(_523_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_405_), .C(_509_), .Y(_524_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_522_), .B(_524_), .Y(_30_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_511_), .C(in125), .Y(_525_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(in125), .Y(_526_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_405_), .C(_514_), .Y(_527_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_525_), .B(_527_), .Y(_31_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_0_), .Y(_528_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_1_), .B(_528_), .Y(_529_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_3_), .Y(_530_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_2_), .B(_530_), .Y(_531_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(out724) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(out725) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(out726) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(out727) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_4_), .Y(out728) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_5_), .Y(out729) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_6_), .Y(out730) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_7_), .Y(out731) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_8_), .Y(out732) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_9_), .Y(out733) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(out734) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(out735) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_12_), .Y(out736) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_13_), .Y(out737) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_14_), .Y(out738) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_15_), .Y(out739) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_16_), .Y(out740) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_17_), .Y(out741) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_18_), .Y(out742) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_19_), .Y(out743) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(out744) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_21_), .Y(out745) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_22_), .Y(out746) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_23_), .Y(out747) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_24_), .Y(out748) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_25_), .Y(out749) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_26_), .Y(out750) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_27_), .Y(out751) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_28_), .Y(out752) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_29_), .Y(out753) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_30_), .Y(out754) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_31_), .Y(out755) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(in69), .B(in65), .Y(_344_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(in69), .B(in65), .Y(_345_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_345_), .Y(_346_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(in73), .B(in77), .Y(_347_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(in73), .B(in77), .Y(_348_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_348_), .B(_347_), .Y(_349_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_349_), .Y(_350_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(in65), .Y(_351_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(in69), .B(_351_), .Y(_352_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(in69), .Y(_353_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(in65), .B(_353_), .Y(_354_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_354_), .Y(_355_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(in73), .Y(_356_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(in77), .B(_356_), .Y(_357_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(in77), .Y(_358_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(in73), .B(_358_), .Y(_359_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_359_), .Y(_360_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_355_), .B(_360_), .Y(_361_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(in17), .B(in1), .Y(_362_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(in33), .B(in49), .Y(_363_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_363_), .B(_362_), .Y(_364_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(in17), .B(in1), .Y(_365_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(in33), .B(in49), .Y(_366_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_366_), .Y(_367_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_367_), .C(_350_), .D(_361_), .Y(_368_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_355_), .Y(_369_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_346_), .B(_360_), .Y(_370_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_366_), .Y(_371_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_363_), .Y(_372_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_372_), .C(_369_), .D(_370_), .Y(_373_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(in129), .B(in137), .Y(_374_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_374_), .Y(_375_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(in85), .B(in81), .Y(_376_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(in85), .B(in81), .Y(_377_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_376_), .B(_377_), .Y(_378_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(in89), .B(in93), .Y(_379_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(in89), .B(in93), .Y(_380_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_380_), .B(_379_), .Y(_381_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_381_), .Y(_382_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(in81), .Y(_383_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(in85), .B(_383_), .Y(_384_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(in85), .Y(_385_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(in81), .B(_385_), .Y(_386_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_386_), .Y(_387_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(in89), .Y(_388_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(in93), .B(_388_), .Y(_389_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(in93), .Y(_390_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(in89), .B(_390_), .Y(_391_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_391_), .Y(_392_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_392_), .Y(_393_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_382_), .C(_375_), .Y(_32_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_387_), .Y(_33_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_392_), .Y(_34_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .C(_374_), .Y(_35_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_32_), .C(_368_), .D(_373_), .Y(_36_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_367_), .C(_369_), .D(_370_), .Y(_37_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_372_), .C(_350_), .D(_361_), .Y(_38_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_382_), .C(_374_), .Y(_39_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .C(_375_), .Y(_40_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_39_), .C(_37_), .D(_38_), .Y(_41_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_41_), .Y(Ckt499b_M1_S_7_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(in101), .B(in97), .Y(_42_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(in105), .B(in109), .Y(_43_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(in105), .B(in109), .Y(_44_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_44_), .C(_42_), .Y(_45_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(in101), .B(in97), .Y(_46_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_43_), .Y(_47_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_46_), .Y(_48_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(in21), .B(in5), .Y(_49_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(in37), .B(in53), .Y(_50_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_50_), .Y(_51_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(in21), .B(in5), .Y(_52_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(in37), .B(in53), .Y(_53_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_52_), .Y(_54_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_48_), .C(_51_), .D(_54_), .Y(_55_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(in105), .B(in109), .Y(_56_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_56_), .Y(_57_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_42_), .Y(_58_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_53_), .Y(_59_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_50_), .Y(_60_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_57_), .C(_59_), .D(_60_), .Y(_61_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(in137), .B(in130), .Y(_62_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(in117), .B(in113), .Y(_63_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(in117), .B(in113), .Y(_64_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(in121), .B(in125), .Y(_65_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(in121), .B(in125), .Y(_66_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_63_), .C(_65_), .D(_66_), .Y(_67_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(in113), .Y(_68_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(in117), .B(_68_), .Y(_69_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(in117), .Y(_70_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(in113), .B(_70_), .Y(_71_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(in121), .Y(_72_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(in125), .B(_72_), .Y(_73_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(in125), .Y(_74_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(in121), .B(_74_), .Y(_75_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_71_), .C(_73_), .D(_75_), .Y(_76_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_76_), .C(_62_), .Y(_77_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_62_), .Y(_78_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .C(_69_), .D(_71_), .Y(_79_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_63_), .C(_73_), .D(_75_), .Y(_80_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_80_), .C(_78_), .Y(_81_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_77_), .Y(_82_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_61_), .C(_82_), .Y(_83_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_46_), .Y(_84_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_56_), .Y(_85_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_52_), .Y(_86_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_50_), .Y(_87_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_84_), .C(_86_), .D(_87_), .Y(_88_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_47_), .B(_42_), .Y(_89_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_56_), .Y(_90_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_50_), .Y(_91_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_53_), .Y(_92_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_89_), .C(_91_), .D(_92_), .Y(_93_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_64_), .Y(_94_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_65_), .Y(_95_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_95_), .Y(_96_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_71_), .Y(_97_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_75_), .Y(_98_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_98_), .Y(_99_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_96_), .C(_62_), .Y(_100_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_97_), .Y(_101_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_98_), .Y(_102_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_102_), .C(_78_), .Y(_103_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_100_), .C(_88_), .D(_93_), .Y(_104_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_83_), .Y(Ckt499b_M1_S_6_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_344_), .C(_347_), .D(_348_), .Y(_105_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_354_), .C(_357_), .D(_359_), .Y(_106_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(in137), .B(in131), .Y(_107_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_106_), .C(_107_), .Y(_108_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_348_), .C(_352_), .D(_354_), .Y(_109_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_344_), .C(_357_), .D(_359_), .Y(_110_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_107_), .Y(_111_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_110_), .C(_111_), .Y(_112_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_108_), .Y(_113_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(in25), .B(in9), .Y(_114_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(in41), .B(in57), .Y(_115_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_115_), .Y(_116_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(in25), .B(in9), .Y(_117_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(in41), .B(in57), .Y(_118_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_117_), .Y(_119_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_48_), .C(_116_), .D(_119_), .Y(_120_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_118_), .Y(_121_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_115_), .Y(_122_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_58_), .B(_57_), .C(_121_), .D(_122_), .Y(_123_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_123_), .C(_113_), .Y(_124_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_350_), .C(_107_), .Y(_125_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_370_), .B(_369_), .C(_111_), .Y(_126_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_117_), .Y(_127_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_115_), .Y(_128_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_84_), .C(_127_), .D(_128_), .Y(_129_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_115_), .Y(_130_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_118_), .Y(_131_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_89_), .C(_130_), .D(_131_), .Y(_132_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_126_), .B(_125_), .C(_129_), .D(_132_), .Y(_133_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_124_), .Y(Ckt499b_M1_S_5_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_376_), .C(_379_), .D(_380_), .Y(_134_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_384_), .B(_386_), .C(_389_), .D(_391_), .Y(_135_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(in137), .B(in132), .Y(_136_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(_136_), .Y(_137_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_380_), .C(_384_), .D(_386_), .Y(_138_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_376_), .C(_389_), .D(_391_), .Y(_139_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_136_), .Y(_140_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .C(_140_), .Y(_141_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_137_), .Y(_142_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(in29), .B(in13), .Y(_143_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(in45), .B(in61), .Y(_144_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_144_), .Y(_145_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(in29), .B(in13), .Y(_146_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(in45), .B(in61), .Y(_147_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_146_), .Y(_148_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_80_), .C(_145_), .D(_148_), .Y(_149_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_147_), .Y(_150_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_144_), .Y(_151_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_76_), .C(_150_), .D(_151_), .Y(_152_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_152_), .C(_142_), .Y(_153_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_382_), .C(_136_), .Y(_154_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .C(_140_), .Y(_155_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_146_), .Y(_156_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_144_), .Y(_157_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .C(_101_), .D(_102_), .Y(_158_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_144_), .Y(_159_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_147_), .Y(_160_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_159_), .B(_160_), .C(_96_), .D(_99_), .Y(_161_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_155_), .B(_154_), .C(_158_), .D(_161_), .Y(_162_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_153_), .Y(Ckt499b_M1_S_4_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(in1), .B(in5), .Y(_163_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(in1), .B(in5), .Y(_164_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_163_), .B(_164_), .Y(_165_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(in9), .B(in13), .Y(_166_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(in9), .B(in13), .Y(_167_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_166_), .Y(_168_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_168_), .Y(_169_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(in5), .Y(_170_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(in1), .B(_170_), .Y(_171_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(in1), .Y(_172_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(in5), .B(_172_), .Y(_173_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_173_), .Y(_174_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(in9), .Y(_175_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(in13), .B(_175_), .Y(_176_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(in13), .Y(_177_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(in9), .B(_177_), .Y(_178_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_178_), .Y(_179_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_179_), .Y(_180_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(in65), .B(in81), .Y(_181_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(in97), .B(in113), .Y(_182_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_181_), .Y(_183_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(in65), .B(in81), .Y(_184_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(in97), .B(in113), .Y(_185_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_185_), .Y(_186_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_186_), .C(_169_), .D(_180_), .Y(_187_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_174_), .Y(_188_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_179_), .Y(_189_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_185_), .Y(_190_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_182_), .Y(_191_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(_188_), .D(_189_), .Y(_192_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(in137), .B(in133), .Y(_193_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_193_), .Y(_194_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(in17), .B(in21), .Y(_195_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(in17), .B(in21), .Y(_196_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_196_), .Y(_197_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(in25), .B(in29), .Y(_198_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(in25), .B(in29), .Y(_199_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_198_), .Y(_200_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_200_), .Y(_201_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(in21), .Y(_202_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(in17), .B(_202_), .Y(_203_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(in17), .Y(_204_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(in21), .B(_204_), .Y(_205_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_205_), .Y(_206_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(in25), .Y(_207_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(in29), .B(_207_), .Y(_208_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(in29), .Y(_209_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(in25), .B(_209_), .Y(_210_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_210_), .Y(_211_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_211_), .Y(_212_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_201_), .C(_194_), .Y(_213_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_200_), .B(_206_), .Y(_214_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_197_), .B(_211_), .Y(_215_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_215_), .C(_193_), .Y(_216_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_216_), .B(_213_), .C(_187_), .D(_192_), .Y(_217_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_186_), .C(_188_), .D(_189_), .Y(_218_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_191_), .C(_169_), .D(_180_), .Y(_219_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_201_), .C(_193_), .Y(_220_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_215_), .C(_194_), .Y(_221_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_220_), .C(_218_), .D(_219_), .Y(_222_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_222_), .Y(Ckt499b_M1_S_3_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(in33), .B(in37), .Y(_223_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(in41), .B(in45), .Y(_224_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(in41), .B(in45), .Y(_225_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .C(_223_), .Y(_226_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(in33), .B(in37), .Y(_227_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_224_), .Y(_228_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_227_), .Y(_229_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(in69), .B(in85), .Y(_230_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(in101), .B(in117), .Y(_231_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .Y(_232_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(in69), .B(in85), .Y(_233_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(in101), .B(in117), .Y(_234_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_233_), .Y(_235_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_229_), .C(_232_), .D(_235_), .Y(_236_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(in41), .B(in45), .Y(_237_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_237_), .Y(_238_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_223_), .Y(_239_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_234_), .Y(_240_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_231_), .Y(_241_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_238_), .C(_240_), .D(_241_), .Y(_242_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(in137), .B(in134), .Y(_243_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(in49), .B(in53), .Y(_244_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(in49), .B(in53), .Y(_245_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(in57), .B(in61), .Y(_246_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(in57), .B(in61), .Y(_247_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_244_), .C(_246_), .D(_247_), .Y(_248_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(in53), .Y(_249_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(in49), .B(_249_), .Y(_250_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(in49), .Y(_251_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(in53), .B(_251_), .Y(_252_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(in57), .Y(_253_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(in61), .B(_253_), .Y(_254_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(in61), .Y(_255_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(in57), .B(_255_), .Y(_256_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_252_), .C(_254_), .D(_256_), .Y(_257_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_257_), .C(_243_), .Y(_258_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_243_), .Y(_259_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_247_), .C(_250_), .D(_252_), .Y(_260_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_245_), .B(_244_), .C(_254_), .D(_256_), .Y(_261_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_261_), .C(_259_), .Y(_262_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_258_), .Y(_263_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_242_), .C(_263_), .Y(_264_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_227_), .Y(_265_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_237_), .Y(_266_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_234_), .B(_233_), .Y(_267_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .Y(_268_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_265_), .C(_267_), .D(_268_), .Y(_269_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_223_), .Y(_270_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_237_), .Y(_271_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_231_), .Y(_272_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_234_), .Y(_273_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_270_), .C(_272_), .D(_273_), .Y(_274_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_245_), .Y(_275_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_246_), .Y(_276_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_276_), .Y(_277_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_252_), .Y(_278_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_256_), .Y(_279_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_279_), .Y(_280_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_280_), .B(_277_), .C(_243_), .Y(_281_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_278_), .Y(_282_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_279_), .Y(_283_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_282_), .B(_283_), .C(_259_), .Y(_284_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_281_), .C(_269_), .D(_274_), .Y(_285_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_264_), .Y(Ckt499b_M1_S_2_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_163_), .C(_166_), .D(_167_), .Y(_286_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_171_), .B(_173_), .C(_176_), .D(_178_), .Y(_287_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(in137), .B(in135), .Y(_288_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_287_), .C(_288_), .Y(_289_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_167_), .C(_171_), .D(_173_), .Y(_290_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_163_), .C(_176_), .D(_178_), .Y(_291_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_288_), .Y(_292_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_290_), .B(_291_), .C(_292_), .Y(_293_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_289_), .Y(_294_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(in73), .B(in89), .Y(_295_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(in105), .B(in121), .Y(_296_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .Y(_297_) );
XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(in73), .B(in89), .Y(_298_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(in105), .B(in121), .Y(_299_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_298_), .Y(_300_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_229_), .C(_297_), .D(_300_), .Y(_301_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_299_), .Y(_302_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_296_), .Y(_303_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_238_), .C(_302_), .D(_303_), .Y(_304_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_304_), .C(_294_), .Y(_305_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_169_), .C(_288_), .Y(_306_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_188_), .C(_292_), .Y(_307_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_298_), .Y(_308_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .Y(_309_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_266_), .B(_265_), .C(_308_), .D(_309_), .Y(_310_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_298_), .B(_296_), .Y(_311_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_299_), .Y(_312_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_270_), .C(_311_), .D(_312_), .Y(_313_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_306_), .C(_310_), .D(_313_), .Y(_314_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_305_), .Y(Ckt499b_M1_S_1_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_195_), .C(_198_), .D(_199_), .Y(_315_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_205_), .C(_208_), .D(_210_), .Y(_316_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(in137), .B(in136), .Y(_317_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_316_), .C(_317_), .Y(_318_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_199_), .C(_203_), .D(_205_), .Y(_319_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_195_), .C(_208_), .D(_210_), .Y(_320_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_317_), .Y(_321_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_320_), .C(_321_), .Y(_322_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_322_), .B(_318_), .Y(_323_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(in77), .B(in93), .Y(_324_) );
XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(in109), .B(in125), .Y(_325_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_325_), .Y(_326_) );
XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(in77), .B(in93), .Y(_327_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(in109), .B(in125), .Y(_328_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_327_), .Y(_329_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_261_), .C(_326_), .D(_329_), .Y(_330_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_328_), .Y(_331_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_325_), .Y(_332_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_257_), .C(_331_), .D(_332_), .Y(_333_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_333_), .C(_323_), .Y(_334_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_201_), .C(_317_), .Y(_335_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_215_), .C(_321_), .Y(_336_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_327_), .Y(_337_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_325_), .Y(_338_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_338_), .C(_282_), .D(_283_), .Y(_339_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_325_), .Y(_340_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_328_), .Y(_341_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_341_), .C(_277_), .D(_280_), .Y(_342_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_335_), .C(_339_), .D(_342_), .Y(_343_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_334_), .Y(Ckt499b_M1_S_0_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_7_), .Y(_532_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_6_), .B(_532_), .Y(_533_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_5_), .B(Ckt499b_M1_S_4_), .Y(_534_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_531_), .C(_533_), .Y(_535_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_535_), .C(in1), .Y(_536_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(in1), .Y(_537_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_1_), .Y(_538_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_0_), .B(_538_), .Y(_539_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_2_), .Y(_540_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_3_), .B(_540_), .Y(_541_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_6_), .Y(_542_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_7_), .B(_542_), .Y(_543_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_5_), .B(Ckt499b_M1_S_4_), .Y(_544_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_541_), .C(_543_), .Y(_545_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_539_), .C(_545_), .Y(_546_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_536_), .B(_546_), .Y(_0_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_7_), .B(_542_), .Y(_547_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_531_), .C(_547_), .Y(_548_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_548_), .C(in5), .Y(_549_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(in5), .Y(_550_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_6_), .B(_532_), .Y(_551_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_541_), .C(_551_), .Y(_552_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_550_), .B(_539_), .C(_552_), .Y(_553_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_553_), .Y(_1_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_5_), .Y(_394_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_4_), .B(_394_), .Y(_395_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_6_), .B(Ckt499b_M1_S_7_), .Y(_396_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_531_), .C(_395_), .Y(_397_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_397_), .C(in9), .Y(_398_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(in9), .Y(_399_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_4_), .Y(_400_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_5_), .B(_400_), .Y(_401_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_6_), .B(Ckt499b_M1_S_7_), .Y(_402_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_541_), .C(_401_), .Y(_403_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_539_), .C(_403_), .Y(_404_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_404_), .Y(_2_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_5_), .B(_400_), .Y(_405_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_531_), .C(_405_), .Y(_406_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_529_), .B(_406_), .C(in13), .Y(_407_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(in13), .Y(_408_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(Ckt499b_M1_S_4_), .B(_394_), .Y(_409_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_541_), .C(_409_), .Y(_410_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_408_), .B(_539_), .C(_410_), .Y(_411_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_407_), .B(_411_), .Y(_3_) );
endmodule
