module o8_cpu ( gnd, vdd, clk_i, rst_i, int_i, data_i, ack_i, err_i, addr_o, data_o, rd_o, wr_o);

input gnd, vdd;
input clk_i;
input rst_i;
input int_i;
input ack_i;
input err_i;
output rd_o;
output wr_o;
input [7:0] data_i;
output [15:0] addr_o;
output [7:0] data_o;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf8) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf7) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf6) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf5) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf4) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf3) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf2) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf1) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk_i), .Y(clk_i_bF_buf0) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf3) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf2) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf1) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_68_), .Y(_68__bF_buf0) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(pg_zf), .Y(pg_zf_bF_buf6) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(pg_zf), .Y(pg_zf_bF_buf5) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(pg_zf), .Y(pg_zf_bF_buf4) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(pg_zf), .Y(pg_zf_bF_buf3) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(pg_zf), .Y(pg_zf_bF_buf2) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(pg_zf), .Y(pg_zf_bF_buf1) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(pg_zf), .Y(pg_zf_bF_buf0) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(autocarry), .B(rst_i), .Y(_10_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(_10_), .Y(_11_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(_12_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(_12_), .Y(_13_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(state_4_), .Y(_14_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_14_), .C(_13_), .Y(_15_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(_16_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(state_0_), .Y(_17_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_14_), .C(_17_), .Y(_18_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_18_), .C(_11_), .Y(ac_sel_0_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(op_cf), .Y(_19_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(ac_sel_0_), .Y(_20_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_20_), .Y(autocarry_next) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf0), .Y(_21_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(state_2_), .C(state_4_), .Y(_22_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_17_), .C(_11_), .Y(_23_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_14_), .Y(_24_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(_25_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_25_), .C(_21_), .Y(_26_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_24_), .Y(_27_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_27_), .Y(_28_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(data_i[0]), .Y(_29_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_25_), .Y(_30_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(_31_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(_32_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_31_), .C(_32_), .Y(_33_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_33_), .C(_18_), .Y(_34_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_10_), .C(_34_), .Y(_35_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(alu_res_0_), .B(ac_sel_0_), .C(_35_), .Y(_36_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_36_), .C(_21_), .Y(_5__0_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(data_i[1]), .Y(_37_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_10_), .C(_34_), .Y(_38_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(alu_res_1_), .B(ac_sel_0_), .C(_38_), .Y(_39_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_39_), .C(_21_), .Y(_5__1_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(data_i[2]), .Y(_40_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_10_), .C(_34_), .Y(_41_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(alu_res_2_), .B(ac_sel_0_), .C(_41_), .Y(_42_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_42_), .C(_21_), .Y(_5__2_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(data_i[3]), .Y(_43_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_10_), .C(_34_), .Y(_44_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(alu_res_3_), .B(ac_sel_0_), .C(_44_), .Y(_45_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_45_), .C(_21_), .Y(_5__3_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(data_i[4]), .Y(_46_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_10_), .C(_34_), .Y(_47_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(alu_res_4_), .B(ac_sel_0_), .C(_47_), .Y(_48_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_48_), .C(_21_), .Y(_5__4_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(data_i[5]), .Y(_49_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_49_), .B(_10_), .C(_34_), .Y(_50_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(alu_res_5_), .B(ac_sel_0_), .C(_50_), .Y(_51_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_51_), .C(_21_), .Y(_5__5_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(data_i[6]), .Y(_52_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_52_), .B(_10_), .C(_34_), .Y(_53_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(alu_res_6_), .B(ac_sel_0_), .C(_53_), .Y(_54_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_54_), .C(_21_), .Y(_5__6_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(data_i[7]), .Y(_55_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_10_), .C(_34_), .Y(_56_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(op_sf), .B(ac_sel_0_), .C(_56_), .Y(_57_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(_57_), .C(_21_), .Y(_5__7_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(state_4_), .C(_16_), .Y(_58_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_22_), .C(_13_), .D(_58_), .Y(_59_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(autocarry), .B(ac_which_2_), .Y(_60_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(autocarry), .B(_59_), .C(_60_), .Y(_61_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(rst_i), .Y(_62_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(autocarry), .B(_18_), .C(_62_), .Y(_63_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_27_), .C(_63_), .Y(_64_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(_64_), .Y(_65_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(autocarry), .Y(_66_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(ac_which_2_), .S(_66_), .Y(_67_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_17_), .C(_22_), .Y(_68_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(pg_zf_bF_buf1), .C(_12_), .Y(_69_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_66_), .B(_22_), .C(_69_), .Y(_70_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_68__bF_buf1), .C(_70_), .Y(_71_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_67_), .C(pg_zf_bF_buf1), .Y(_72_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_36_), .B(_65_), .C(_72_), .Y(_1__8_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_65_), .C(_72_), .Y(_1__9_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_65_), .C(_72_), .Y(_1__10_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_65_), .C(_72_), .Y(_1__11_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_65_), .C(_72_), .Y(_1__12_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_65_), .C(_72_), .Y(_1__13_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_54_), .B(_65_), .C(_72_), .Y(_1__14_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_65_), .C(_72_), .Y(_1__15_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_18_), .C(pg_zf_bF_buf1), .Y(_73_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(_36_), .C(_73_), .Y(_2__0_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(_39_), .C(_73_), .Y(_2__1_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(_42_), .C(_73_), .Y(_2__2_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(_45_), .C(_73_), .Y(_2__3_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf3), .B(_48_), .C(_73_), .Y(_2__4_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf2), .B(_51_), .C(_73_), .Y(_2__5_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf1), .B(_54_), .C(_73_), .Y(_2__6_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_68__bF_buf0), .B(_57_), .C(_73_), .Y(_2__7_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(autocarry), .B(_62_), .Y(_74_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_74_), .C(_68__bF_buf1), .Y(_9__0_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_74_), .Y(_9__1_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_74_), .Y(_9__2_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_74_), .Y(_9__3_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_74_), .Y(_9__4_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(prev_cf), .Y(_75_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_74_), .C(_20_), .Y(alu_cf) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(rst_i), .B(_21_), .Y(_76_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_76_), .Y(_77_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_27_), .B(_34_), .C(_66_), .Y(_78_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_60_), .C(_77_), .Y(_7__7_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_78_), .Y(_4__7_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(alu_res_0_), .Y(_79_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_68__bF_buf0), .C(_73_), .Y(_1__0_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(alu_res_1_), .Y(_80_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_80_), .B(_68__bF_buf2), .C(_73_), .Y(_1__1_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(alu_res_2_), .Y(_81_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_81_), .B(_68__bF_buf2), .C(_73_), .Y(_1__2_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(alu_res_3_), .Y(_82_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_68__bF_buf3), .C(_73_), .Y(_1__3_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(alu_res_4_), .Y(_83_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_68__bF_buf3), .C(_73_), .Y(_1__4_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(alu_res_5_), .Y(_84_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_68__bF_buf3), .C(_73_), .Y(_1__5_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(alu_res_6_), .Y(_85_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_68__bF_buf1), .C(_73_), .Y(_1__6_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(op_sf), .Y(_86_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_68__bF_buf0), .C(_73_), .Y(_1__7_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(op_zf), .Y(_87_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_28_), .C(_21_), .Y(_0__0_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_28_), .C(_21_), .Y(_0__1_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(alu_of_out), .Y(_88_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_28_), .C(_21_), .Y(_0__2_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(op_sf), .Y(_89_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_28_), .C(_21_), .Y(_0__3_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(op_sf), .Y(_90_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_28_), .C(_21_), .Y(_0__4_) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(ac_sel_0_), .Y(_93_) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf0), .Y(_6__0_) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf3), .Y(_6__1_) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf5), .Y(_6__2_) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf5), .Y(_6__3_) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf3), .Y(_6__4_) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf6), .Y(_6__5_) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf0), .Y(_6__6_) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf6), .Y(_6__7_) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf6), .Y(_3__0_) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf2), .Y(_3__1_) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf6), .Y(_3__2_) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf1), .Y(_3__3_) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf4), .Y(_3__4_) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf6), .Y(_3__5_) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf6), .Y(_3__6_) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf4), .Y(_3__7_) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf3), .Y(_3__8_) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf5), .Y(_3__9_) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf2), .Y(_3__10_) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf5), .Y(_3__11_) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf0), .Y(_3__12_) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf4), .Y(_3__13_) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf5), .Y(_3__14_) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf2), .Y(_3__15_) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf3), .Y(_8__0_) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf2), .Y(_8__1_) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf0), .Y(_8__2_) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf2), .Y(_8__3_) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf4), .Y(_8__4_) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf5), .Y(_8__5_) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf2), .Y(_8__6_) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf3), .Y(_8__7_) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf5), .Y(_8__8_) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf1), .Y(_8__9_) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf6), .Y(_8__10_) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf0), .Y(_8__11_) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf4), .Y(_8__12_) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf1), .Y(_8__13_) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf3), .Y(_8__14_) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf4), .Y(_8__15_) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf4), .Y(_0__5_) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[0]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[1]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[2]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[3]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[4]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[5]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[6]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(addr_o[7]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[8]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[9]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[10]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[11]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[12]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[13]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[14]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(addr_o[15]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[0]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[1]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[2]) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[3]) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[4]) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[5]) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[6]) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(_92__7_), .Y(data_o[7]) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(rd_o) );
BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(wr_o) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(ac_sel_0_), .Q(ac_which_2_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_5__0_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_5__1_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(_5__2_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_5__3_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_5__4_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_5__5_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(_5__6_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_5__7_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_6__0_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_6__1_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_6__2_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_6__3_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_6__4_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_6__5_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_6__6_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_6__7_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_3__0_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_3__1_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_3__2_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_3__3_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_3__4_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_3__5_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_3__6_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_3__7_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_3__8_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_3__9_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_3__10_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_3__11_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_3__12_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_3__13_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_3__14_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_3__15_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_8__0_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_8__1_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_8__2_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_8__3_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_8__4_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_8__5_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_8__6_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_8__7_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_8__8_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_8__9_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_8__10_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf1), .D(_8__11_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_8__12_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_8__13_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_8__14_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(_8__15_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_0__0_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(_0__1_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_0__2_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_0__3_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_0__4_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf0), .D(_0__5_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_1__0_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_1__1_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(_1__2_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_1__3_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_1__4_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_1__5_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_1__6_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_1__7_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_1__8_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_1__9_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_1__10_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_1__11_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_1__12_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_1__13_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_1__14_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_1__15_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_2__0_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_2__1_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf5), .D(_2__2_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf6), .D(_2__3_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf3), .D(_2__4_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf8), .D(_2__5_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_2__6_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf4), .D(_2__7_), .Q(pg_zf) );
DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(_9__0_), .Q(state_0_) );
DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(_9__1_), .Q(state_1_) );
DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_9__2_), .Q(state_2_) );
DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_9__3_), .Q(state_3_) );
DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf7), .D(_9__4_), .Q(state_4_) );
DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(op_cf), .Q(prev_cf) );
DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_i_bF_buf2), .D(autocarry_next), .Q(autocarry) );
$_DLATCH_P_ $_DLATCH_P__1 ( .gnd(gnd), .vdd(vdd), .D(gnd), .E(rst_i), .Q(pg_zf) );
$_DLATCH_P_ $_DLATCH_P__2 ( .gnd(gnd), .vdd(vdd), .D(pg_zf), .E(vdd), .Q(_92__7_) );
$_DLATCH_P_ $_DLATCH_P__3 ( .gnd(gnd), .vdd(vdd), .D(_4__7_), .E(vdd), .Q(_91__7_) );
$_DLATCH_P_ $_DLATCH_P__4 ( .gnd(gnd), .vdd(vdd), .D(_7__7_), .E(vdd), .Q(_91__15_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(alu_rsx_7_), .B(gnd), .Y(op_sf) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(alu_rsx_6_), .Y(alu_res_6_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(alu_rsx_5_), .Y(alu_res_5_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(alu_rsx_4_), .Y(alu_res_4_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(alu_rsx_3_), .Y(alu_res_3_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(alu_rsx_2_), .Y(alu_res_2_) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(alu_rsx_1_), .Y(_285_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_285_), .Y(alu_res_1_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(alu_rsx_0_), .Y(_286_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_286_), .Y(alu_res_0_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(alu_res_3_), .B(alu_res_2_), .Y(_287_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_286_), .C(_287_), .Y(_288_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(op_sf), .B(alu_res_6_), .Y(_289_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(alu_res_5_), .B(alu_res_4_), .Y(_290_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_290_), .Y(_291_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_288_), .Y(op_zf) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .B(_91__15_), .Y(_292_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(op_sf), .Y(_293_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .B(_91__15_), .Y(_294_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(op_sf), .B(_294_), .C(_293_), .Y(alu_of_out) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_295_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf3), .B(_295_), .Y(_296_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_296_), .Y(_297_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_297_), .Y(_299_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(_299_), .Y(_300_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(alu_cf), .Y(_301_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(_302_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_302_), .Y(_303_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_304_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .B(_304_), .Y(_305_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_306_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .B(_306_), .Y(_307_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(_308_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_308_), .Y(_309_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_305_), .C(_307_), .D(_309_), .Y(_310_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_311_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_312_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_313_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_314_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_312_), .C(_313_), .D(_314_), .Y(_315_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_310_), .Y(_316_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_316_), .B(_301_), .Y(_317_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(pg_zf_bF_buf2), .Y(_319_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_319_), .Y(_320_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .B(_304_), .Y(_321_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_302_), .Y(_322_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_308_), .Y(_323_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .B(_306_), .Y(_324_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_321_), .B(_322_), .C(_323_), .D(_324_), .Y(_95_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(_96_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf1), .B(_96_), .Y(_97_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_97_), .Y(_98_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(pg_zf_bF_buf0), .B(_295_), .Y(_99_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_99_), .Y(_100_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_101_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_102_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_101_), .Y(_103_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_103_), .Y(_104_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_98_), .C(_100_), .D(_104_), .Y(_105_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_316_), .C(_105_), .Y(_106_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_108_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_109_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_108_), .Y(_110_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(pg_zf_bF_buf6), .Y(_111_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_111_), .Y(_325_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_325_), .Y(_112_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_319_), .B(_112_), .C(_320_), .Y(_113_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_97_), .Y(_114_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_307_), .B(_309_), .C(_114_), .Y(_115_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_113_), .C(_115_), .Y(_116_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_106_), .Y(_117_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_317_), .C(_117_), .Y(_298_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .Y(_118_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_118_), .Y(_119_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .B(_304_), .Y(_120_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .Y(_121_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_121_), .Y(_122_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .B(_306_), .Y(_123_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_119_), .B(_120_), .C(_122_), .D(_123_), .Y(_125_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_121_), .Y(_126_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_127_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_102_), .C(_126_), .D(_127_), .Y(_128_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_125_), .Y(_129_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_129_), .Y(_130_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(alu_cf), .B(_315_), .C(_95_), .Y(_131_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_131_), .C(_300_), .Y(_132_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_130_), .B(_131_), .C(_132_), .Y(_133_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_110_), .C(_103_), .Y(_134_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_297_), .Y(_135_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_305_), .C(alu_cf), .Y(_136_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(_136_), .Y(_137_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_137_), .Y(_138_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(_138_), .Y(_139_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(_320_), .Y(_140_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_141_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_125_), .Y(_142_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_123_), .Y(_143_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_144_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_143_), .C(_100_), .D(_144_), .Y(_145_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_142_), .C(_145_), .Y(_146_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_129_), .C(_146_), .Y(_147_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_139_), .Y(_148_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_133_), .Y(_149_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_103_), .C(_149_), .Y(_318_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_150_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_151_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .Y(_152_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_153_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_144_), .Y(_154_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_308_), .Y(_155_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_156_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_109_), .C(_155_), .D(_156_), .Y(_157_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_301_), .B(_157_), .C(_310_), .Y(_158_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_129_), .C(_125_), .Y(_159_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_154_), .C(_159_), .Y(_160_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_154_), .Y(_161_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_131_), .C(_142_), .Y(_162_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_161_), .B(_162_), .C(_299_), .Y(_163_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_137_), .Y(_164_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(_135_), .Y(_165_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_150_), .C(_165_), .Y(_166_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_161_), .Y(_167_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_153_), .Y(_168_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_169_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_169_), .C(_98_), .D(_168_), .Y(_170_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_171_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_151_), .C(_144_), .D(_171_), .Y(_172_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_170_), .B(_167_), .C(_172_), .Y(_173_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_166_), .C(_173_), .Y(_174_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_163_), .C(_174_), .Y(_107_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_175_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_175_), .Y(_176_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_177_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_178_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_178_), .Y(_179_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_176_), .Y(_180_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_168_), .B(_160_), .Y(_181_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_180_), .Y(_182_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_180_), .B(_181_), .C(_299_), .Y(_183_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_169_), .C(_137_), .Y(_184_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_164_), .B(_177_), .C(_165_), .Y(_185_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_141_), .Y(_186_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_187_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(_188_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_175_), .C(_100_), .D(_188_), .Y(_189_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_113_), .C(_189_), .Y(_190_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_190_), .Y(_191_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_180_), .C(_191_), .Y(_192_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_185_), .C(_192_), .Y(_193_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_183_), .C(_193_), .Y(_124_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_194_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(_194_), .Y(_195_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_195_), .Y(_196_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_187_), .B(_194_), .Y(_197_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_197_), .Y(_198_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(_198_), .Y(_199_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_154_), .C(_180_), .Y(_200_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_153_), .C(_176_), .Y(_201_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_201_), .C(_162_), .D(_200_), .Y(_202_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_202_), .Y(_203_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_176_), .B(_179_), .C(_161_), .Y(_204_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_175_), .C(_201_), .Y(_205_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_159_), .C(_205_), .Y(_206_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_206_), .C(_299_), .Y(_207_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_187_), .Y(_208_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_187_), .C(_165_), .Y(_209_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_196_), .Y(_210_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_211_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(_211_), .Y(_212_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_114_), .C(_100_), .D(_212_), .Y(_213_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_187_), .C(_213_), .Y(_214_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_210_), .C(_214_), .Y(_215_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_199_), .C(_215_), .Y(_216_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_209_), .C(_216_), .Y(_217_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_207_), .C(_217_), .Y(_94__4_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_218_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_218_), .Y(_219_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_212_), .Y(_220_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_218_), .Y(_221_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_221_), .Y(_222_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_202_), .C(_196_), .Y(_223_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_222_), .Y(_224_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_223_), .C(_299_), .Y(_225_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_212_), .Y(_226_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_226_), .Y(_227_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_211_), .C(_165_), .Y(_228_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__7_), .Y(_229_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_229_), .Y(_230_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_114_), .C(_100_), .D(_230_), .Y(_231_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_220_), .C(_231_), .Y(_232_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_140_), .C(_232_), .Y(_233_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_211_), .C(_233_), .Y(_234_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_227_), .C(_234_), .Y(_235_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .C(_235_), .Y(_94__5_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(_91__15_), .Y(_236_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_230_), .Y(_237_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_236_), .Y(_238_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_238_), .Y(_239_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(_239_), .Y(_240_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_222_), .Y(_241_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_218_), .C(_196_), .Y(_242_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_212_), .B(_219_), .C(_242_), .Y(_243_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_202_), .C(_243_), .Y(_244_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_240_), .C(_300_), .Y(_245_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_244_), .C(_245_), .Y(_246_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_229_), .C(_165_), .Y(_247_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_229_), .C(_247_), .Y(_248_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_237_), .Y(_249_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_91__7_), .B(gnd), .Y(_250_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(_250_), .Y(_251_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_251_), .C(_98_), .D(_249_), .Y(_252_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_239_), .C(_252_), .Y(_253_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_236_), .B(_114_), .Y(_254_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_113_), .C(_254_), .Y(_255_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_253_), .Y(_256_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_256_), .C(_246_), .Y(_94__6_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_244_), .Y(_257_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_91__15_), .B(gnd), .Y(_258_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_258_), .Y(_259_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_258_), .Y(_260_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_259_), .Y(_261_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_261_), .Y(_262_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_262_), .Y(_263_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_257_), .C(_263_), .Y(_264_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_222_), .Y(_265_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_242_), .C(_265_), .D(_206_), .Y(_266_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_261_), .Y(_267_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_249_), .B(_267_), .Y(_268_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_266_), .C(_268_), .Y(_269_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_299_), .B(_269_), .Y(_270_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_229_), .C(_184_), .Y(_271_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_251_), .C(_165_), .Y(_272_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_271_), .B(_251_), .C(_272_), .Y(_273_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_258_), .Y(_274_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_251_), .C(_274_), .Y(_275_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_113_), .C(_275_), .Y(_276_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_140_), .C(_276_), .Y(_277_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_273_), .B(_277_), .Y(_278_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_264_), .B(_270_), .C(_278_), .Y(_94__7_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_259_), .Y(_279_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_240_), .Y(_280_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_280_), .C(_279_), .Y(_281_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_280_), .Y(_282_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_206_), .B(_282_), .C(_281_), .Y(_283_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_135_), .B(_251_), .C(_271_), .Y(_284_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_283_), .C(_284_), .Y(_94__8_) );
$_DLATCH_P_ $_DLATCH_P__5 ( .gnd(gnd), .vdd(vdd), .D(_298_), .E(_325_), .Q(alu_rsx_0_) );
$_DLATCH_P_ $_DLATCH_P__6 ( .gnd(gnd), .vdd(vdd), .D(_318_), .E(_325_), .Q(alu_rsx_1_) );
$_DLATCH_P_ $_DLATCH_P__7 ( .gnd(gnd), .vdd(vdd), .D(_107_), .E(_325_), .Q(alu_rsx_2_) );
$_DLATCH_P_ $_DLATCH_P__8 ( .gnd(gnd), .vdd(vdd), .D(_124_), .E(_325_), .Q(alu_rsx_3_) );
$_DLATCH_P_ $_DLATCH_P__9 ( .gnd(gnd), .vdd(vdd), .D(_94__4_), .E(_325_), .Q(alu_rsx_4_) );
$_DLATCH_P_ $_DLATCH_P__10 ( .gnd(gnd), .vdd(vdd), .D(_94__5_), .E(_325_), .Q(alu_rsx_5_) );
$_DLATCH_P_ $_DLATCH_P__11 ( .gnd(gnd), .vdd(vdd), .D(_94__6_), .E(_325_), .Q(alu_rsx_6_) );
