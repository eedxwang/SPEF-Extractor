module rle_enc ( gnd, vdd, clk, rst, recv_ready, send_ready, in_data, end_of_stream, rd_req, out_data, wr_req);

input gnd, vdd;
input clk;
input rst;
input recv_ready;
input send_ready;
input end_of_stream;
output rd_req;
output wr_req;
input [7:0] in_data;
output [23:0] out_data;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf3) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf2) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf1) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(state_7_), .Y(state_7_bF_buf0) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(_7_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(state_8_), .Y(_8_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(end_of_stream), .Y(_9_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .C(_7_), .Y(_206__0_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .B(_7_), .Y(_10_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(recv_ready), .Y(_11_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_207__3_), .Y(_12_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_207__2_), .Y(_13_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .B(_207__0_), .Y(_14_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .C(_14_), .Y(_15_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(_207__7_), .Y(_16_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_207__6_), .Y(_17_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_207__5_), .B(_207__4_), .Y(_18_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .C(_18_), .Y(_19_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_19_), .Y(_20_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_207__16_), .Y(_21_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_207__19_), .Y(_22_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_207__18_), .Y(_23_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_22_), .C(_23_), .Y(_24_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_207__20_), .Y(_25_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_207__17_), .Y(_26_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_207__22_), .B(_207__21_), .Y(_27_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_26_), .C(_27_), .Y(_28_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_28_), .Y(_29_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_207__9_), .Y(_30_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_207__8_), .Y(_31_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_207__11_), .B(_207__10_), .Y(_32_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_31_), .C(_32_), .Y(_33_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_207__15_), .Y(_34_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(_207__14_), .Y(_35_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_207__13_), .B(_207__12_), .Y(_36_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_35_), .C(_36_), .Y(_37_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_37_), .Y(_38_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_38_), .B(_29_), .Y(_39_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_20_), .C(_9_), .Y(_40_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(shift_count_1_), .B(shift_count_0_), .C(shift_count_2_), .Y(_41_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(shift_count_3_), .B(_41_), .Y(_42_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(_43_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(new_bitstream), .B(_43_), .Y(_44_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_44_), .Y(_45_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_45_), .C(_7_), .Y(_46_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_40_), .C(_46_), .Y(_206__5_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_47_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(new_bitstream), .Y(_48_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_43_), .Y(_49_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(state_6_), .Y(_50_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(send_ready), .B(_50_), .Y(_51_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_51_), .B(_49_), .C(_7_), .Y(_52_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_11_), .B(_47_), .C(_52_), .Y(_206__6_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(shift_count_3_), .B(_41_), .C(_44_), .Y(_53_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(state_8_), .C(state_1_), .Y(_54_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_53_), .B(_54_), .C(rst), .Y(_206__7_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(shift_count_0_), .B(_44_), .Y(_55_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(state_5_), .Y(_56_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_43_), .C(_49_), .Y(_57_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(shift_count_0_), .C(_55_), .Y(_4__0_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(shift_count_0_), .Y(_58_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(new_bitstream), .B(_58_), .Y(_59_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(shift_count_1_), .B(_59_), .Y(_60_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_60_), .Y(_61_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_61_), .Y(_62_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(state_2_), .C(_62_), .Y(_63_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(state_2_), .C(shift_count_1_), .Y(_64_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_63_), .Y(_4__1_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_62_), .S(shift_count_2_), .Y(_4__2_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_61_), .B(shift_count_2_), .Y(_65_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_45_), .Y(_66_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_56_), .C(shift_count_3_), .Y(_67_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_65_), .C(_66_), .Y(_4__3_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_0_), .Y(_68_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(_69_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(state_1_), .Y(_70_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_70_), .Y(_71_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_43_), .C(_71_), .Y(_72_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_72_), .Y(_73_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[0]), .C(shift_buf_1_), .D(_44_), .Y(_74_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_73_), .C(_74_), .Y(_3__0_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_1_), .B(_72_), .Y(_75_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[1]), .Y(_76_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_2_), .B(_44_), .Y(_77_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_76_), .B(_77_), .C(_75_), .Y(_3__1_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_2_), .B(_72_), .Y(_78_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[2]), .Y(_79_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_3_), .B(_44_), .Y(_80_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_80_), .C(_78_), .Y(_3__2_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_3_), .B(_72_), .Y(_81_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[3]), .Y(_82_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_4_), .B(_44_), .Y(_83_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_83_), .C(_81_), .Y(_3__3_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_4_), .B(_72_), .Y(_84_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[4]), .Y(_85_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_5_), .B(_44_), .Y(_86_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_86_), .C(_84_), .Y(_3__4_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_5_), .B(_72_), .Y(_87_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[5]), .Y(_88_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_6_), .B(_44_), .Y(_89_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_89_), .C(_87_), .Y(_3__5_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_6_), .B(_72_), .Y(_90_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[6]), .Y(_91_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_7_), .B(_44_), .Y(_92_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_91_), .B(_92_), .C(_90_), .Y(_3__6_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_7_), .Y(_93_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .B(in_data[7]), .Y(_94_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_93_), .B(_73_), .C(_94_), .Y(_3__7_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_0_), .B(value_type), .C(new_bitstream), .Y(_95_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_0_), .B(value_type), .C(_95_), .Y(_96_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(state_7_bF_buf2), .Y(_97_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf2), .Y(_98_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_98_), .Y(_99_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_97_), .C(_99_), .D(_96_), .Y(_1_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(new_bitstream), .B(state_7_bF_buf2), .Y(_100_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_98_), .C(value_type), .Y(_101_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_68_), .B(_100_), .C(_101_), .Y(_5_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_69_), .Y(_102_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_102_), .C(_56_), .Y(_2_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_209_), .B(_69_), .Y(_103_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_103_), .C(_50_), .Y(_6_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_207__0_), .B(_96_), .Y(_104_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_97_), .Y(_105_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(_105_), .Y(_106_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_207__0_), .Y(_107_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(shift_buf_0_), .B(value_type), .Y(_108_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_95_), .C(_107_), .Y(_109_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_109_), .Y(_110_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_207__0_), .B(_106_), .C(state_7_bF_buf1), .D(_110_), .Y(_111_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_111_), .Y(_0__0_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .Y(_112_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_207__1_), .C(_98_), .Y(_113_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .B(_109_), .C(_113_), .Y(_114_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_105_), .C(_114_), .Y(_0__1_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_112_), .B(_110_), .C(_13_), .Y(_115_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .B(_207__2_), .C(_109_), .Y(_116_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(_116_), .C(_115_), .Y(_117_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_105_), .C(_117_), .Y(_0__2_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_116_), .B(_12_), .Y(_118_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(state_7_bF_buf1), .C(_106_), .Y(_119_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_116_), .C(_12_), .Y(_120_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_120_), .Y(_121_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_119_), .Y(_0__3_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_207__4_), .Y(_122_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(_122_), .Y(_123_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_118_), .B(_123_), .C(_122_), .D(_119_), .Y(_0__4_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_207__5_), .Y(_124_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .B(_207__2_), .Y(_125_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_207__4_), .B(_207__0_), .C(_207__3_), .Y(_126_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_126_), .Y(_127_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_127_), .B(_96_), .Y(_128_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_207__5_), .C(_98_), .Y(_129_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_207__5_), .B(_128_), .C(_129_), .Y(_130_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_105_), .C(_130_), .Y(_0__5_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_96_), .B(_127_), .Y(_131_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_131_), .C(_17_), .Y(_132_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_207__5_), .B(_207__6_), .C(_128_), .Y(_133_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf1), .B(_132_), .C(_133_), .Y(_134_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_17_), .B(_105_), .C(_134_), .Y(_0__6_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_207__7_), .B(_106_), .Y(_135_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_133_), .C(state_7_bF_buf1), .Y(_136_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_133_), .C(_135_), .D(_136_), .Y(_0__7_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_133_), .C(_31_), .Y(_137_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_207__5_), .B(_207__7_), .Y(_138_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_207__6_), .B(_207__8_), .Y(_139_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_138_), .B(_139_), .Y(_140_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_96_), .C(_127_), .Y(_141_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf0), .B(_141_), .C(_137_), .Y(_142_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_31_), .B(_105_), .C(_142_), .Y(_0__8_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_207__9_), .B(_140_), .Y(_143_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_143_), .Y(_144_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_207__9_), .B(_106_), .C(state_7_bF_buf0), .D(_144_), .Y(_145_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_141_), .C(_145_), .Y(_0__9_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_207__10_), .Y(_146_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_131_), .Y(_147_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_147_), .B(_207__10_), .C(_98_), .Y(_148_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_207__10_), .B(_147_), .C(_148_), .Y(_149_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_105_), .C(_149_), .Y(_0__10_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_106_), .B(_148_), .C(_207__11_), .Y(_150_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_207__10_), .B(state_7_bF_buf0), .C(_147_), .Y(_151_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_207__11_), .B(_151_), .C(_150_), .Y(_0__11_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_207__12_), .Y(_152_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_207__11_), .B(_207__10_), .Y(_153_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_144_), .C(_152_), .Y(_154_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_153_), .Y(_155_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_207__12_), .B(_155_), .C(_147_), .Y(_156_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf0), .B(_156_), .C(_154_), .Y(_157_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_152_), .B(_105_), .C(_157_), .Y(_0__12_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_207__13_), .Y(_158_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(_207__13_), .B(_106_), .Y(_159_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_30_), .B(_141_), .Y(_160_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_207__13_), .B(_207__12_), .Y(_161_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_161_), .Y(_162_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_160_), .Y(_163_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf3), .B(_163_), .Y(_164_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_156_), .C(_159_), .D(_164_), .Y(_0__13_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_207__14_), .B(_106_), .Y(_165_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_163_), .C(state_7_bF_buf0), .Y(_166_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_35_), .B(_163_), .C(_165_), .D(_166_), .Y(_0__14_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_207__14_), .B(_162_), .C(_160_), .Y(_167_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_207__15_), .B(_106_), .Y(_168_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_35_), .Y(_169_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_169_), .C(_160_), .Y(_170_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf3), .B(_170_), .Y(_171_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_34_), .B(_167_), .C(_168_), .D(_171_), .Y(_0__15_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_207__16_), .B(_106_), .Y(_172_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_207__15_), .B(_207__14_), .C(_207__16_), .Y(_173_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_163_), .C(state_7_bF_buf3), .Y(_174_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_170_), .C(_172_), .D(_174_), .Y(_0__16_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_173_), .Y(_175_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_175_), .C(_160_), .Y(_176_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_207__17_), .B(_106_), .Y(_177_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_173_), .Y(_178_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_178_), .Y(_179_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_163_), .C(state_7_bF_buf3), .Y(_180_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_26_), .B(_176_), .C(_177_), .D(_180_), .Y(_0__17_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_178_), .C(_160_), .Y(_181_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_207__18_), .B(_106_), .Y(_182_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_207__18_), .B(_178_), .Y(_183_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_183_), .B(_163_), .C(state_7_bF_buf3), .Y(_184_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_181_), .C(_182_), .D(_184_), .Y(_0__18_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_183_), .Y(_185_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_185_), .C(_160_), .Y(_186_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_207__19_), .B(_106_), .Y(_187_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_207__19_), .B(_207__18_), .C(_178_), .Y(_188_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_163_), .C(state_7_bF_buf3), .Y(_189_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_186_), .C(_187_), .D(_189_), .Y(_0__19_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_163_), .C(_25_), .Y(_190_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_207__9_), .B(_207__20_), .C(_162_), .Y(_191_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_188_), .C(_141_), .Y(_192_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_25_), .B(_105_), .C(_98_), .D(_192_), .Y(_193_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_193_), .Y(_0__20_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_188_), .Y(_194_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_191_), .B(_141_), .Y(_195_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_207__21_), .B(_194_), .C(_195_), .Y(_196_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_97_), .C(state_7_bF_buf2), .D(_196_), .Y(_197_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_192_), .B(state_7_bF_buf2), .C(_207__21_), .Y(_198_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_197_), .Y(_0__21_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_207__22_), .Y(_199_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(state_7_bF_buf2), .B(_199_), .Y(_200_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_200_), .Y(_201_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_197_), .C(_201_), .Y(_0__22_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(state_3_), .Y(_204_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(send_ready), .B(_7_), .Y(_202_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_202_), .Y(_205_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(recv_ready), .Y(_203_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_10_), .Y(_206__3_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(rst), .B(_98_), .Y(_206__2_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_7_), .B(state_4_), .Y(_206__8_) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_207__0_), .Y(out_data[0]) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_207__1_), .Y(out_data[1]) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_207__2_), .Y(out_data[2]) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_207__3_), .Y(out_data[3]) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_207__4_), .Y(out_data[4]) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_207__5_), .Y(out_data[5]) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_207__6_), .Y(out_data[6]) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_207__7_), .Y(out_data[7]) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_207__8_), .Y(out_data[8]) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_207__9_), .Y(out_data[9]) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_207__10_), .Y(out_data[10]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_207__11_), .Y(out_data[11]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_207__12_), .Y(out_data[12]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_207__13_), .Y(out_data[13]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_207__14_), .Y(out_data[14]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_207__15_), .Y(out_data[15]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_207__16_), .Y(out_data[16]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_207__17_), .Y(out_data[17]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_207__18_), .Y(out_data[18]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_207__19_), .Y(out_data[19]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_207__20_), .Y(out_data[20]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_207__21_), .Y(out_data[21]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_207__22_), .Y(out_data[22]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(value_type), .Y(out_data[23]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_208_), .Y(rd_req) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_209_), .Y(wr_req) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_206__0_), .Q(state_0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_204_), .Q(state_1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_206__2_), .Q(state_2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_206__3_), .Q(state_3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_205_), .Q(state_4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_206__5_), .Q(state_5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_206__6_), .Q(state_6_) );
DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_206__7_), .Q(state_7_) );
DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_206__8_), .Q(state_8_) );
DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_2_), .Q(_208_) );
DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_6_), .Q(_209_) );
DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__0_), .Q(_207__0_) );
DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__1_), .Q(_207__1_) );
DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__2_), .Q(_207__2_) );
DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__3_), .Q(_207__3_) );
DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__4_), .Q(_207__4_) );
DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__5_), .Q(_207__5_) );
DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__6_), .Q(_207__6_) );
DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__7_), .Q(_207__7_) );
DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__8_), .Q(_207__8_) );
DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__9_), .Q(_207__9_) );
DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__10_), .Q(_207__10_) );
DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__11_), .Q(_207__11_) );
DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__12_), .Q(_207__12_) );
DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__13_), .Q(_207__13_) );
DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__14_), .Q(_207__14_) );
DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__15_), .Q(_207__15_) );
DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__16_), .Q(_207__16_) );
DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__17_), .Q(_207__17_) );
DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__18_), .Q(_207__18_) );
DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__19_), .Q(_207__19_) );
DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__20_), .Q(_207__20_) );
DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__21_), .Q(_207__21_) );
DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__22_), .Q(_207__22_) );
DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4__0_), .Q(shift_count_0_) );
DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4__1_), .Q(shift_count_1_) );
DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4__2_), .Q(shift_count_2_) );
DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_4__3_), .Q(shift_count_3_) );
DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_5_), .Q(value_type) );
DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3__0_), .Q(shift_buf_0_) );
DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3__1_), .Q(shift_buf_1_) );
DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3__2_), .Q(shift_buf_2_) );
DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3__3_), .Q(shift_buf_3_) );
DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3__4_), .Q(shift_buf_4_) );
DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3__5_), .Q(shift_buf_5_) );
DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3__6_), .Q(shift_buf_6_) );
DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3__7_), .Q(shift_buf_7_) );
DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_1_), .Q(new_bitstream) );
endmodule
