module spi_master ( gnd, vdd, clk, rst, data_in, MISO, send, MOSI, SCLK, SS, done);

input gnd, vdd;
input clk;
input rst;
input MISO;
input send;
output MOSI;
output SCLK;
output SS;
output done;
input [6:0] data_in;

NAND2X1 NAND2X1_1 (  .A(load), .B(data_in[3]), .Y(_41_) );
OAI21X1 OAI21X1_1 (  .A(load), .B(_40_), .C(_41_), .Y(_27_) );
MUX2X1 MUX2X1_1 (  .A(shift_data[3]), .B(shift_data[4]), .S(shift_en), .Y(_42_) );
NAND2X1 NAND2X1_2 (  .A(load), .B(data_in[4]), .Y(_43_) );
OAI21X1 OAI21X1_2 (  .A(load), .B(_42_), .C(_43_), .Y(_28_) );
MUX2X1 MUX2X1_2 (  .A(shift_data[4]), .B(shift_data[5]), .S(shift_en), .Y(_44_) );
NAND2X1 NAND2X1_3 (  .A(load), .B(data_in[5]), .Y(_45_) );
OAI21X1 OAI21X1_3 (  .A(load), .B(_44_), .C(_45_), .Y(_29_) );
MUX2X1 MUX2X1_3 (  .A(shift_data[5]), .B(shift_data[6]), .S(shift_en), .Y(_46_) );
NAND2X1 NAND2X1_4 (  .A(load), .B(data_in[6]), .Y(_47_) );
OAI21X1 OAI21X1_4 (  .A(load), .B(_46_), .C(_47_), .Y(_30_) );
MUX2X1 MUX2X1_4 (  .A(shift_data[6]), .B(_0_), .S(shift_en), .Y(_48_) );
NOR2X1 NOR2X1_1 (  .A(load), .B(_48_), .Y(_33_) );
INVX2 INVX2_1 (  .A(clk), .Y(_36_) );
INVX4 INVX4_1 (  .A(rst), .Y(_38_) );
DFFSR DFFSR_1 (  .CLK(_36_), .D(_49_), .Q(shift_data[0]), .R(_38_), .S(vdd) );
DFFSR DFFSR_2 (  .CLK(_36_), .D(_25_), .Q(shift_data[1]), .R(_38_), .S(vdd) );
DFFSR DFFSR_3 (  .CLK(_36_), .D(_26_), .Q(shift_data[2]), .R(_38_), .S(vdd) );
DFFSR DFFSR_4 (  .CLK(_36_), .D(_27_), .Q(shift_data[3]), .R(_38_), .S(vdd) );
DFFSR DFFSR_5 (  .CLK(_36_), .D(_28_), .Q(shift_data[4]), .R(_38_), .S(vdd) );
DFFSR DFFSR_6 (  .CLK(_36_), .D(_29_), .Q(shift_data[5]), .R(_38_), .S(vdd) );
DFFSR DFFSR_7 (  .CLK(_36_), .D(_30_), .Q(shift_data[6]), .R(_38_), .S(vdd) );
DFFSR DFFSR_8 (  .CLK(_36_), .D(_33_), .Q(_0_), .R(_38_), .S(vdd) );
BUFX2 BUFX2_1 (  .A(_0_), .Y(MOSI) );
BUFX2 BUFX2_2 (  .A(_1_), .Y(SCLK) );
BUFX2 BUFX2_3 (  .A(_2_), .Y(SS) );
BUFX2 BUFX2_4 (  .A(_3_), .Y(done) );
INVX1 INVX1_1 (  .A(ctrl_cstate[1]), .Y(_5_) );
NAND3X1 NAND3X1_1 (  .A(ctrl_count[0]), .B(ctrl_count[1]), .C(ctrl_count[2]), .Y(_6_) );
NAND2X1 NAND2X1_5 (  .A(ctrl_clk_en), .B(_6_), .Y(_7_) );
NAND2X1 NAND2X1_6 (  .A(_5_), .B(_7_), .Y(_22_) );
INVX1 INVX1_2 (  .A(ctrl_clk_en), .Y(_8_) );
INVX1 INVX1_3 (  .A(ctrl_cstate[4]), .Y(_9_) );
OAI22X1 OAI22X1_1 (  .A(_9_), .B(send), .C(_8_), .D(_6_), .Y(_23_[4]) );
NAND2X1 NAND2X1_7 (  .A(ctrl_clk_en), .B(ctrl_count[0]), .Y(_4_[0]) );
NAND2X1 NAND2X1_8 (  .A(ctrl_count[0]), .B(ctrl_count[1]), .Y(_11_) );
INVX1 INVX1_4 (  .A(_11_), .Y(_13_) );
NOR2X1 NOR2X1_2 (  .A(ctrl_count[0]), .B(ctrl_count[1]), .Y(_15_) );
OAI21X1 OAI21X1_5 (  .A(_15_), .B(_13_), .C(ctrl_clk_en), .Y(_4_[1]) );
NAND2X1 NAND2X1_9 (  .A(ctrl_count[2]), .B(_11_), .Y(_16_) );
INVX1 INVX1_5 (  .A(ctrl_count[2]), .Y(_17_) );
NAND3X1 NAND3X1_2 (  .A(ctrl_count[0]), .B(ctrl_count[1]), .C(_17_), .Y(_18_) );
NAND3X1 NAND3X1_3 (  .A(ctrl_clk_en), .B(_18_), .C(_16_), .Y(_4_[2]) );
NOR2X1 NOR2X1_3 (  .A(ctrl_cstate[4]), .B(ctrl_cstate[3]), .Y(_19_) );
OAI21X1 OAI21X1_6 (  .A(ctrl_cstate[1]), .B(ctrl_clk_en), .C(_19_), .Y(_2_) );
INVX1 INVX1_6 (  .A(clk), .Y(_14_) );
NOR2X1 NOR2X1_4 (  .A(_8_), .B(_14_), .Y(_1_) );
OAI21X1 OAI21X1_7 (  .A(ctrl_cstate[4]), .B(ctrl_cstate[0]), .C(send), .Y(_20_) );
INVX1 INVX1_7 (  .A(_20_), .Y(_10_) );
INVX1 INVX1_8 (  .A(ctrl_cstate[0]), .Y(_21_) );
NOR2X1 NOR2X1_5 (  .A(send), .B(_21_), .Y(_12_) );
INVX4 INVX4_2 (  .A(rst), .Y(_24_) );
BUFX2 BUFX2_5 (  .A(ctrl_cstate[4]), .Y(_3_) );
BUFX4 BUFX4_1 (  .A(ctrl_cstate[3]), .Y(load) );
BUFX4 BUFX4_2 (  .A(ctrl_clk_en), .Y(shift_en) );
DFFSR DFFSR_9 (  .CLK(clk), .D(_12_), .Q(ctrl_cstate[0]), .R(vdd), .S(_24_) );
DFFSR DFFSR_10 (  .CLK(clk), .D(ctrl_cstate[3]), .Q(ctrl_cstate[1]), .R(_24_), .S(vdd) );
DFFSR DFFSR_11 (  .CLK(clk), .D(_22_), .Q(ctrl_clk_en), .R(_24_), .S(vdd) );
DFFSR DFFSR_12 (  .CLK(clk), .D(_10_), .Q(ctrl_cstate[3]), .R(_24_), .S(vdd) );
DFFSR DFFSR_13 (  .CLK(clk), .D(_23_[4]), .Q(ctrl_cstate[4]), .R(_24_), .S(vdd) );
DFFSR DFFSR_14 (  .CLK(_14_), .D(_4_[0]), .Q(ctrl_count[0]), .R(vdd), .S(_24_) );
DFFSR DFFSR_15 (  .CLK(_14_), .D(_4_[1]), .Q(ctrl_count[1]), .R(vdd), .S(_24_) );
DFFSR DFFSR_16 (  .CLK(_14_), .D(_4_[2]), .Q(ctrl_count[2]), .R(vdd), .S(_24_) );
MUX2X1 MUX2X1_5 (  .A(MISO), .B(shift_data[0]), .S(shift_en), .Y(_31_) );
NAND2X1 NAND2X1_10 (  .A(data_in[0]), .B(load), .Y(_32_) );
OAI21X1 OAI21X1_8 (  .A(load), .B(_31_), .C(_32_), .Y(_49_) );
MUX2X1 MUX2X1_6 (  .A(shift_data[0]), .B(shift_data[1]), .S(shift_en), .Y(_34_) );
NAND2X1 NAND2X1_11 (  .A(load), .B(data_in[1]), .Y(_35_) );
OAI21X1 OAI21X1_9 (  .A(load), .B(_34_), .C(_35_), .Y(_25_) );
MUX2X1 MUX2X1_7 (  .A(shift_data[1]), .B(shift_data[2]), .S(shift_en), .Y(_37_) );
NAND2X1 NAND2X1_12 (  .A(load), .B(data_in[2]), .Y(_39_) );
OAI21X1 OAI21X1_10 (  .A(load), .B(_37_), .C(_39_), .Y(_26_) );
MUX2X1 MUX2X1_8 (  .A(shift_data[2]), .B(shift_data[3]), .S(shift_en), .Y(_40_) );
endmodule
