module spi_master ( gnd, vdd, clk, rst, data_in, MISO, send, MOSI, SCLK, SS, done);

input gnd, vdd;
input clk;
input rst;
input MISO;
input send;
output MOSI;
output SCLK;
output SS;
output done;
input [6:0] data_in;

NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(load), .B(data_in[3]), .Y(_41_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_40_), .C(_41_), .Y(_27_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(shift_data_3_), .B(shift_data_4_), .S(shift_en), .Y(_42_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(load), .B(data_in[4]), .Y(_43_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_42_), .C(_43_), .Y(_28_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(shift_data_4_), .B(shift_data_5_), .S(shift_en), .Y(_44_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(load), .B(data_in[5]), .Y(_45_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_44_), .C(_45_), .Y(_29_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(shift_data_5_), .B(shift_data_6_), .S(shift_en), .Y(_46_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(load), .B(data_in[6]), .Y(_47_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_46_), .C(_47_), .Y(_30_) );
MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(shift_data_6_), .B(_0_), .S(shift_en), .Y(_48_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_48_), .Y(_33_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(_36_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(_38_) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_49_), .Q(shift_data_0_), .R(_38_), .S(vdd) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_25_), .Q(shift_data_1_), .R(_38_), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_26_), .Q(shift_data_2_), .R(_38_), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_27_), .Q(shift_data_3_), .R(_38_), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_28_), .Q(shift_data_4_), .R(_38_), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_29_), .Q(shift_data_5_), .R(_38_), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_30_), .Q(shift_data_6_), .R(_38_), .S(vdd) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(_36_), .D(_33_), .Q(_0_), .R(_38_), .S(vdd) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_0_), .Y(MOSI) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_1_), .Y(SCLK) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_2_), .Y(SS) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_3_), .Y(done) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_1_), .Y(_5_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(ctrl_count_0_), .B(ctrl_count_1_), .C(ctrl_count_2_), .Y(_6_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(ctrl_clk_en), .B(_6_), .Y(_7_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_5_), .B(_7_), .Y(_22_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(ctrl_clk_en), .Y(_8_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_4_), .Y(_9_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_9_), .B(send), .C(_8_), .D(_6_), .Y(_23__4_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(ctrl_clk_en), .B(ctrl_count_0_), .Y(_4__0_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(ctrl_count_0_), .B(ctrl_count_1_), .Y(_11_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_11_), .Y(_13_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(ctrl_count_0_), .B(ctrl_count_1_), .Y(_15_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_15_), .B(_13_), .C(ctrl_clk_en), .Y(_4__1_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(ctrl_count_2_), .B(_11_), .Y(_16_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(ctrl_count_2_), .Y(_17_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(ctrl_count_0_), .B(ctrl_count_1_), .C(_17_), .Y(_18_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(ctrl_clk_en), .B(_18_), .C(_16_), .Y(_4__2_) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_4_), .B(ctrl_cstate_3_), .Y(_19_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_1_), .B(ctrl_clk_en), .C(_19_), .Y(_2_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(_14_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_14_), .Y(_1_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_4_), .B(ctrl_cstate_0_), .C(send), .Y(_20_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_20_), .Y(_10_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_0_), .Y(_21_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(send), .B(_21_), .Y(_12_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(rst), .Y(_24_) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_4_), .Y(_3_) );
BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(ctrl_cstate_3_), .Y(load) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(ctrl_clk_en), .Y(shift_en) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_12_), .Q(ctrl_cstate_0_), .R(vdd), .S(_24_) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(ctrl_cstate_3_), .Q(ctrl_cstate_1_), .R(_24_), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_22_), .Q(ctrl_clk_en), .R(_24_), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_10_), .Q(ctrl_cstate_3_), .R(_24_), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(_23__4_), .Q(ctrl_cstate_4_), .R(_24_), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_4__0_), .Q(ctrl_count_0_), .R(vdd), .S(_24_) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_4__1_), .Q(ctrl_count_1_), .R(vdd), .S(_24_) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(_14_), .D(_4__2_), .Q(ctrl_count_2_), .R(vdd), .S(_24_) );
MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(MISO), .B(shift_data_0_), .S(shift_en), .Y(_31_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(data_in[0]), .B(load), .Y(_32_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_31_), .C(_32_), .Y(_49_) );
MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(shift_data_0_), .B(shift_data_1_), .S(shift_en), .Y(_34_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(load), .B(data_in[1]), .Y(_35_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_34_), .C(_35_), .Y(_25_) );
MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(shift_data_1_), .B(shift_data_2_), .S(shift_en), .Y(_37_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(load), .B(data_in[2]), .Y(_39_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(load), .B(_37_), .C(_39_), .Y(_26_) );
MUX2X1 MUX2X1_8 ( .gnd(gnd), .vdd(vdd), .A(shift_data_2_), .B(shift_data_3_), .S(shift_en), .Y(_40_) );
endmodule
